module moduleName #(
    parameter DATA_WIDTH = 32;
) (
    ports
);
    
endmodule